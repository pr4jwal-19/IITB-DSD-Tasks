library ieee;
use ieee.std_logic_1164.all;

library work;
use work.Gates.all;

entity FourBitAdder_1 is
 
	PORT (a0,a1,a2,a3,b0,b1,b2,b3,cin1: in std_logic;  s0,s1,s2,s3,cout:out std_logic);

end entity;

architecture halfadder of FourBitAdder_1 is 
	signal sig1,sig2,sig3,sig4,sig5,sig6,sig7:std_logic;
begin 
      inst1: XOR_2 port map(A => b0,B =>cin1,Y => sig1);
		inst2: XOR_2 port map(A => b1,B =>cin1,Y => sig2);
		inst3: XOR_2 port map(A => b2,B =>cin1,Y => sig3);
		inst4: XOR_2 port map(A => b3,B =>cin1,Y => sig4);
      inst5: FULL_ADDER port map(A => a0,B =>sig1,CIN =>cin1,S=>s0,C => sig5);
		inst6: FULL_ADDER port map(A => a1,B =>sig2,CIN => sig5,S=>s1,C=> sig6);
		inst7: FULL_ADDER port map(A => a2,B =>sig3,CIN => sig6,S=>s2,C=> sig7);
		inst8: FULL_ADDER port map(A => a3,B =>sig4,CIN => sig7,S=>s3,C=> cout);

end architecture ;